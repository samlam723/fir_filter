
module dff_16bit_0 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_14 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_13 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_12 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_11 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_10 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_9 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_8 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_7 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_6 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_5 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_4 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_3 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_2 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module dff_16bit_1 ( d, clk, reset, q );
  input [15:0] d;
  output [15:0] q;
  input clk, reset;


  DFFR_X1 q_reg_15_ ( .D(d[15]), .CK(clk), .RN(reset), .Q(q[15]) );
  DFFR_X1 q_reg_14_ ( .D(d[14]), .CK(clk), .RN(reset), .Q(q[14]) );
  DFFR_X1 q_reg_13_ ( .D(d[13]), .CK(clk), .RN(reset), .Q(q[13]) );
  DFFR_X1 q_reg_12_ ( .D(d[12]), .CK(clk), .RN(reset), .Q(q[12]) );
  DFFR_X1 q_reg_11_ ( .D(d[11]), .CK(clk), .RN(reset), .Q(q[11]) );
  DFFR_X1 q_reg_10_ ( .D(d[10]), .CK(clk), .RN(reset), .Q(q[10]) );
  DFFR_X1 q_reg_9_ ( .D(d[9]), .CK(clk), .RN(reset), .Q(q[9]) );
  DFFR_X1 q_reg_8_ ( .D(d[8]), .CK(clk), .RN(reset), .Q(q[8]) );
  DFFR_X1 q_reg_7_ ( .D(d[7]), .CK(clk), .RN(reset), .Q(q[7]) );
  DFFR_X1 q_reg_6_ ( .D(d[6]), .CK(clk), .RN(reset), .Q(q[6]) );
  DFFR_X1 q_reg_5_ ( .D(d[5]), .CK(clk), .RN(reset), .Q(q[5]) );
  DFFR_X1 q_reg_4_ ( .D(d[4]), .CK(clk), .RN(reset), .Q(q[4]) );
  DFFR_X1 q_reg_3_ ( .D(d[3]), .CK(clk), .RN(reset), .Q(q[3]) );
  DFFR_X1 q_reg_2_ ( .D(d[2]), .CK(clk), .RN(reset), .Q(q[2]) );
  DFFR_X1 q_reg_1_ ( .D(d[1]), .CK(clk), .RN(reset), .Q(q[1]) );
  DFFR_X1 q_reg_0_ ( .D(d[0]), .CK(clk), .RN(reset), .Q(q[0]) );
endmodule


module fir_16tap_DW_mult_uns_10 ( a, b, product );
  input [15:0] a;
  input [3:0] b;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  HA_X1 U2 ( .A(a[15]), .B(n2), .CO(product[19]), .S(product[18]) );
  FA_X1 U3 ( .A(a[15]), .B(a[14]), .CI(n3), .CO(n2), .S(product[17]) );
  FA_X1 U4 ( .A(a[14]), .B(a[13]), .CI(n4), .CO(n3), .S(product[16]) );
  FA_X1 U5 ( .A(a[13]), .B(a[12]), .CI(n5), .CO(n4), .S(product[15]) );
  FA_X1 U6 ( .A(a[12]), .B(a[11]), .CI(n6), .CO(n5), .S(product[14]) );
  FA_X1 U7 ( .A(a[11]), .B(a[10]), .CI(n7), .CO(n6), .S(product[13]) );
  FA_X1 U8 ( .A(a[10]), .B(a[9]), .CI(n8), .CO(n7), .S(product[12]) );
  FA_X1 U9 ( .A(a[9]), .B(a[8]), .CI(n9), .CO(n8), .S(product[11]) );
  FA_X1 U10 ( .A(a[8]), .B(a[7]), .CI(n10), .CO(n9), .S(product[10]) );
  FA_X1 U11 ( .A(a[7]), .B(a[6]), .CI(n11), .CO(n10), .S(product[9]) );
  FA_X1 U12 ( .A(a[6]), .B(a[5]), .CI(n12), .CO(n11), .S(product[8]) );
  FA_X1 U13 ( .A(a[5]), .B(a[4]), .CI(n13), .CO(n12), .S(product[7]) );
  FA_X1 U14 ( .A(a[4]), .B(a[3]), .CI(n14), .CO(n13), .S(product[6]) );
  FA_X1 U15 ( .A(a[3]), .B(a[2]), .CI(n15), .CO(n14), .S(product[5]) );
  FA_X1 U16 ( .A(a[2]), .B(a[1]), .CI(n16), .CO(n15), .S(product[4]) );
  HA_X1 U17 ( .A(a[0]), .B(a[1]), .CO(n16), .S(product[3]) );
  CLKBUF_X1 U22 ( .A(a[0]), .Z(product[2]) );
endmodule


module fir_16tap_DW_mult_uns_9 ( a, b, product );
  input [15:0] a;
  input [3:0] b;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  HA_X1 U2 ( .A(a[15]), .B(n2), .CO(product[19]), .S(product[18]) );
  HA_X1 U3 ( .A(a[14]), .B(n3), .CO(n2), .S(product[17]) );
  HA_X1 U4 ( .A(a[13]), .B(n4), .CO(n3), .S(product[16]) );
  FA_X1 U5 ( .A(a[15]), .B(a[12]), .CI(n5), .CO(n4), .S(product[15]) );
  FA_X1 U6 ( .A(a[14]), .B(a[11]), .CI(n6), .CO(n5), .S(product[14]) );
  FA_X1 U7 ( .A(a[13]), .B(a[10]), .CI(n7), .CO(n6), .S(product[13]) );
  FA_X1 U8 ( .A(a[12]), .B(a[9]), .CI(n8), .CO(n7), .S(product[12]) );
  FA_X1 U9 ( .A(a[11]), .B(a[8]), .CI(n9), .CO(n8), .S(product[11]) );
  FA_X1 U10 ( .A(a[10]), .B(a[7]), .CI(n10), .CO(n9), .S(product[10]) );
  FA_X1 U11 ( .A(a[9]), .B(a[6]), .CI(n11), .CO(n10), .S(product[9]) );
  FA_X1 U12 ( .A(a[8]), .B(a[5]), .CI(n12), .CO(n11), .S(product[8]) );
  FA_X1 U13 ( .A(a[7]), .B(a[4]), .CI(n13), .CO(n12), .S(product[7]) );
  FA_X1 U14 ( .A(a[6]), .B(a[3]), .CI(n14), .CO(n13), .S(product[6]) );
  FA_X1 U15 ( .A(a[5]), .B(a[2]), .CI(n15), .CO(n14), .S(product[5]) );
  FA_X1 U16 ( .A(a[4]), .B(a[1]), .CI(n16), .CO(n15), .S(product[4]) );
  HA_X1 U17 ( .A(a[0]), .B(a[3]), .CO(n16), .S(product[3]) );
  CLKBUF_X1 U22 ( .A(a[2]), .Z(product[2]) );
  CLKBUF_X1 U23 ( .A(a[1]), .Z(product[1]) );
  CLKBUF_X1 U24 ( .A(a[0]), .Z(product[0]) );
endmodule


module fir_16tap_DW_mult_uns_8 ( a, b, product );
  input [15:0] a;
  input [1:0] b;
  output [17:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  HA_X1 U2 ( .A(a[15]), .B(n2), .CO(product[17]), .S(product[16]) );
  FA_X1 U3 ( .A(a[15]), .B(a[14]), .CI(n3), .CO(n2), .S(product[15]) );
  FA_X1 U4 ( .A(a[14]), .B(a[13]), .CI(n4), .CO(n3), .S(product[14]) );
  FA_X1 U5 ( .A(a[13]), .B(a[12]), .CI(n5), .CO(n4), .S(product[13]) );
  FA_X1 U6 ( .A(a[12]), .B(a[11]), .CI(n6), .CO(n5), .S(product[12]) );
  FA_X1 U7 ( .A(a[11]), .B(a[10]), .CI(n7), .CO(n6), .S(product[11]) );
  FA_X1 U8 ( .A(a[10]), .B(a[9]), .CI(n8), .CO(n7), .S(product[10]) );
  FA_X1 U9 ( .A(a[9]), .B(a[8]), .CI(n9), .CO(n8), .S(product[9]) );
  FA_X1 U10 ( .A(a[8]), .B(a[7]), .CI(n10), .CO(n9), .S(product[8]) );
  FA_X1 U11 ( .A(a[7]), .B(a[6]), .CI(n11), .CO(n10), .S(product[7]) );
  FA_X1 U12 ( .A(a[6]), .B(a[5]), .CI(n12), .CO(n11), .S(product[6]) );
  FA_X1 U13 ( .A(a[5]), .B(a[4]), .CI(n13), .CO(n12), .S(product[5]) );
  FA_X1 U14 ( .A(a[4]), .B(a[3]), .CI(n14), .CO(n13), .S(product[4]) );
  FA_X1 U15 ( .A(a[3]), .B(a[2]), .CI(n15), .CO(n14), .S(product[3]) );
  FA_X1 U16 ( .A(a[2]), .B(a[1]), .CI(n16), .CO(n15), .S(product[2]) );
  HA_X1 U17 ( .A(a[0]), .B(a[1]), .CO(n16), .S(product[1]) );
  CLKBUF_X1 U21 ( .A(a[0]), .Z(product[0]) );
endmodule


module fir_16tap_DW_mult_uns_7 ( a, b, product );
  input [15:0] a;
  input [2:0] b;
  output [18:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  HA_X1 U2 ( .A(a[15]), .B(n2), .CO(product[18]), .S(product[17]) );
  FA_X1 U3 ( .A(a[15]), .B(a[14]), .CI(n3), .CO(n2), .S(product[16]) );
  FA_X1 U4 ( .A(a[14]), .B(a[13]), .CI(n4), .CO(n3), .S(product[15]) );
  FA_X1 U5 ( .A(a[13]), .B(a[12]), .CI(n5), .CO(n4), .S(product[14]) );
  FA_X1 U6 ( .A(a[12]), .B(a[11]), .CI(n6), .CO(n5), .S(product[13]) );
  FA_X1 U7 ( .A(a[11]), .B(a[10]), .CI(n7), .CO(n6), .S(product[12]) );
  FA_X1 U8 ( .A(a[10]), .B(a[9]), .CI(n8), .CO(n7), .S(product[11]) );
  FA_X1 U9 ( .A(a[9]), .B(a[8]), .CI(n9), .CO(n8), .S(product[10]) );
  FA_X1 U10 ( .A(a[8]), .B(a[7]), .CI(n10), .CO(n9), .S(product[9]) );
  FA_X1 U11 ( .A(a[7]), .B(a[6]), .CI(n11), .CO(n10), .S(product[8]) );
  FA_X1 U12 ( .A(a[6]), .B(a[5]), .CI(n12), .CO(n11), .S(product[7]) );
  FA_X1 U13 ( .A(a[5]), .B(a[4]), .CI(n13), .CO(n12), .S(product[6]) );
  FA_X1 U14 ( .A(a[4]), .B(a[3]), .CI(n14), .CO(n13), .S(product[5]) );
  FA_X1 U15 ( .A(a[3]), .B(a[2]), .CI(n15), .CO(n14), .S(product[4]) );
  FA_X1 U16 ( .A(a[2]), .B(a[1]), .CI(n16), .CO(n15), .S(product[3]) );
  HA_X1 U17 ( .A(a[0]), .B(a[1]), .CO(n16), .S(product[2]) );
  CLKBUF_X1 U22 ( .A(a[0]), .Z(product[1]) );
endmodule


module fir_16tap_DW01_add_12 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [20:2] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  AND2_X1 U2 ( .A1(A[20]), .A2(carry[20]), .ZN(SUM[21]) );
  XOR2_X1 U3 ( .A(A[20]), .B(carry[20]), .Z(SUM[20]) );
  XOR2_X1 U4 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fir_16tap_DW_mult_uns_6 ( a, b, product );
  input [15:0] a;
  input [2:0] b;
  output [18:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95;

  FA_X1 U6 ( .A(a[12]), .B(n78), .CI(n4), .CO(n3), .S(product[15]) );
  FA_X1 U7 ( .A(a[11]), .B(n79), .CI(n5), .CO(n4), .S(product[14]) );
  FA_X1 U8 ( .A(a[10]), .B(n80), .CI(n6), .CO(n5), .S(product[13]) );
  FA_X1 U9 ( .A(a[9]), .B(n81), .CI(n7), .CO(n6), .S(product[12]) );
  FA_X1 U10 ( .A(a[8]), .B(n82), .CI(n8), .CO(n7), .S(product[11]) );
  FA_X1 U11 ( .A(a[7]), .B(n83), .CI(n9), .CO(n8), .S(product[10]) );
  FA_X1 U12 ( .A(a[6]), .B(n84), .CI(n10), .CO(n9), .S(product[9]) );
  FA_X1 U13 ( .A(a[5]), .B(n85), .CI(n11), .CO(n10), .S(product[8]) );
  FA_X1 U14 ( .A(a[4]), .B(n86), .CI(n12), .CO(n11), .S(product[7]) );
  FA_X1 U15 ( .A(a[3]), .B(n87), .CI(n13), .CO(n12), .S(product[6]) );
  FA_X1 U16 ( .A(a[2]), .B(n88), .CI(n14), .CO(n13), .S(product[5]) );
  FA_X1 U17 ( .A(a[1]), .B(n89), .CI(n15), .CO(n14), .S(product[4]) );
  FA_X1 U18 ( .A(a[0]), .B(n90), .CI(n16), .CO(n15), .S(product[3]) );
  HA_X1 U19 ( .A(n91), .B(n17), .CO(n16), .S(product[2]) );
  HA_X1 U20 ( .A(n92), .B(n93), .CO(n17), .S(product[1]) );
  INV_X1 U41 ( .A(a[1]), .ZN(n92) );
  INV_X1 U42 ( .A(a[0]), .ZN(n93) );
  INV_X1 U43 ( .A(a[15]), .ZN(n78) );
  INV_X1 U44 ( .A(a[3]), .ZN(n90) );
  INV_X1 U45 ( .A(a[4]), .ZN(n89) );
  INV_X1 U46 ( .A(a[5]), .ZN(n88) );
  INV_X1 U47 ( .A(a[6]), .ZN(n87) );
  INV_X1 U48 ( .A(a[7]), .ZN(n86) );
  INV_X1 U49 ( .A(a[8]), .ZN(n85) );
  INV_X1 U50 ( .A(a[9]), .ZN(n84) );
  INV_X1 U51 ( .A(a[10]), .ZN(n83) );
  INV_X1 U52 ( .A(a[11]), .ZN(n82) );
  INV_X1 U53 ( .A(a[12]), .ZN(n81) );
  INV_X1 U54 ( .A(a[13]), .ZN(n80) );
  INV_X1 U55 ( .A(a[2]), .ZN(n91) );
  INV_X1 U56 ( .A(a[14]), .ZN(n79) );
  CLKBUF_X1 U57 ( .A(a[0]), .Z(product[0]) );
  XNOR2_X1 U58 ( .A(a[15]), .B(n94), .ZN(product[18]) );
  NAND2_X1 U59 ( .A1(n95), .A2(n79), .ZN(n94) );
  XNOR2_X1 U60 ( .A(n79), .B(n95), .ZN(product[17]) );
  NOR2_X1 U61 ( .A1(n3), .A2(a[13]), .ZN(n95) );
  XNOR2_X1 U62 ( .A(a[13]), .B(n3), .ZN(product[16]) );
endmodule


module fir_16tap_DW_mult_uns_5 ( a, b, product );
  input [15:0] a;
  input [2:0] b;
  output [18:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  HA_X1 U2 ( .A(a[15]), .B(n2), .CO(product[18]), .S(product[17]) );
  HA_X1 U3 ( .A(a[14]), .B(n3), .CO(n2), .S(product[16]) );
  FA_X1 U4 ( .A(a[15]), .B(a[13]), .CI(n4), .CO(n3), .S(product[15]) );
  FA_X1 U5 ( .A(a[14]), .B(a[12]), .CI(n5), .CO(n4), .S(product[14]) );
  FA_X1 U6 ( .A(a[13]), .B(a[11]), .CI(n6), .CO(n5), .S(product[13]) );
  FA_X1 U7 ( .A(a[12]), .B(a[10]), .CI(n7), .CO(n6), .S(product[12]) );
  FA_X1 U8 ( .A(a[11]), .B(a[9]), .CI(n8), .CO(n7), .S(product[11]) );
  FA_X1 U9 ( .A(a[10]), .B(a[8]), .CI(n9), .CO(n8), .S(product[10]) );
  FA_X1 U10 ( .A(a[9]), .B(a[7]), .CI(n10), .CO(n9), .S(product[9]) );
  FA_X1 U11 ( .A(a[8]), .B(a[6]), .CI(n11), .CO(n10), .S(product[8]) );
  FA_X1 U12 ( .A(a[7]), .B(a[5]), .CI(n12), .CO(n11), .S(product[7]) );
  FA_X1 U13 ( .A(a[6]), .B(a[4]), .CI(n13), .CO(n12), .S(product[6]) );
  FA_X1 U14 ( .A(a[5]), .B(a[3]), .CI(n14), .CO(n13), .S(product[5]) );
  FA_X1 U15 ( .A(a[4]), .B(a[2]), .CI(n15), .CO(n14), .S(product[4]) );
  FA_X1 U16 ( .A(a[3]), .B(a[1]), .CI(n16), .CO(n15), .S(product[3]) );
  HA_X1 U17 ( .A(a[0]), .B(a[2]), .CO(n16), .S(product[2]) );
  CLKBUF_X1 U22 ( .A(a[1]), .Z(product[1]) );
  CLKBUF_X1 U23 ( .A(a[0]), .Z(product[0]) );
endmodule


module fir_16tap_DW01_add_11 ( A, B, CI, SUM, CO );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [18:2] carry;

  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(SUM[19]), .S(SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module fir_16tap_DW_mult_uns_4 ( a, b, product );
  input [15:0] a;
  input [3:0] b;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  FA_X1 U2 ( .A(n18), .B(a[15]), .CI(n2), .CO(product[19]), .S(product[18]) );
  FA_X1 U3 ( .A(n19), .B(n20), .CI(n3), .CO(n2), .S(product[17]) );
  FA_X1 U4 ( .A(n22), .B(n21), .CI(n4), .CO(n3), .S(product[16]) );
  FA_X1 U5 ( .A(n23), .B(n24), .CI(n5), .CO(n4), .S(product[15]) );
  FA_X1 U6 ( .A(n25), .B(n26), .CI(n6), .CO(n5), .S(product[14]) );
  FA_X1 U7 ( .A(n27), .B(n28), .CI(n7), .CO(n6), .S(product[13]) );
  FA_X1 U8 ( .A(n29), .B(n30), .CI(n8), .CO(n7), .S(product[12]) );
  FA_X1 U9 ( .A(n31), .B(n32), .CI(n9), .CO(n8), .S(product[11]) );
  FA_X1 U10 ( .A(n33), .B(n34), .CI(n10), .CO(n9), .S(product[10]) );
  FA_X1 U11 ( .A(n35), .B(n36), .CI(n11), .CO(n10), .S(product[9]) );
  FA_X1 U12 ( .A(n37), .B(n38), .CI(n12), .CO(n11), .S(product[8]) );
  FA_X1 U13 ( .A(n39), .B(n40), .CI(n13), .CO(n12), .S(product[7]) );
  FA_X1 U14 ( .A(n41), .B(n42), .CI(n14), .CO(n13), .S(product[6]) );
  FA_X1 U15 ( .A(n43), .B(n44), .CI(n15), .CO(n14), .S(product[5]) );
  FA_X1 U16 ( .A(n45), .B(n46), .CI(n16), .CO(n15), .S(product[4]) );
  FA_X1 U17 ( .A(n17), .B(a[0]), .CI(n47), .CO(n16), .S(product[3]) );
  HA_X1 U18 ( .A(a[0]), .B(a[2]), .CO(n17), .S(product[2]) );
  HA_X1 U19 ( .A(a[15]), .B(a[14]), .CO(n18), .S(n19) );
  HA_X1 U20 ( .A(a[14]), .B(a[13]), .CO(n20), .S(n21) );
  FA_X1 U21 ( .A(a[12]), .B(a[15]), .CI(a[13]), .CO(n22), .S(n23) );
  FA_X1 U22 ( .A(a[11]), .B(a[14]), .CI(a[12]), .CO(n24), .S(n25) );
  FA_X1 U23 ( .A(a[10]), .B(a[13]), .CI(a[11]), .CO(n26), .S(n27) );
  FA_X1 U24 ( .A(a[9]), .B(a[12]), .CI(a[10]), .CO(n28), .S(n29) );
  FA_X1 U25 ( .A(a[8]), .B(a[11]), .CI(a[9]), .CO(n30), .S(n31) );
  FA_X1 U26 ( .A(a[7]), .B(a[10]), .CI(a[8]), .CO(n32), .S(n33) );
  FA_X1 U27 ( .A(a[6]), .B(a[9]), .CI(a[7]), .CO(n34), .S(n35) );
  FA_X1 U28 ( .A(a[5]), .B(a[8]), .CI(a[6]), .CO(n36), .S(n37) );
  FA_X1 U29 ( .A(a[4]), .B(a[7]), .CI(a[5]), .CO(n38), .S(n39) );
  FA_X1 U30 ( .A(a[3]), .B(a[6]), .CI(a[4]), .CO(n40), .S(n41) );
  FA_X1 U31 ( .A(a[2]), .B(a[5]), .CI(a[3]), .CO(n42), .S(n43) );
  FA_X1 U32 ( .A(a[1]), .B(a[4]), .CI(a[2]), .CO(n44), .S(n45) );
  HA_X1 U33 ( .A(a[3]), .B(a[1]), .CO(n46), .S(n47) );
  CLKBUF_X1 U38 ( .A(a[1]), .Z(product[1]) );
  CLKBUF_X1 U39 ( .A(a[0]), .Z(product[0]) );
endmodule


module fir_16tap_DW_mult_uns_3 ( a, b, product );
  input [15:0] a;
  input [3:0] b;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;

  HA_X1 U2 ( .A(a[15]), .B(n2), .CO(product[19]), .S(product[18]) );
  HA_X1 U3 ( .A(a[14]), .B(n3), .CO(n2), .S(product[17]) );
  FA_X1 U4 ( .A(a[15]), .B(a[13]), .CI(n4), .CO(n3), .S(product[16]) );
  FA_X1 U5 ( .A(a[14]), .B(a[12]), .CI(n5), .CO(n4), .S(product[15]) );
  FA_X1 U6 ( .A(a[13]), .B(a[11]), .CI(n6), .CO(n5), .S(product[14]) );
  FA_X1 U7 ( .A(a[12]), .B(a[10]), .CI(n7), .CO(n6), .S(product[13]) );
  FA_X1 U8 ( .A(a[11]), .B(a[9]), .CI(n8), .CO(n7), .S(product[12]) );
  FA_X1 U9 ( .A(a[10]), .B(a[8]), .CI(n9), .CO(n8), .S(product[11]) );
  FA_X1 U10 ( .A(a[9]), .B(a[7]), .CI(n10), .CO(n9), .S(product[10]) );
  FA_X1 U11 ( .A(a[8]), .B(a[6]), .CI(n11), .CO(n10), .S(product[9]) );
  FA_X1 U12 ( .A(a[7]), .B(a[5]), .CI(n12), .CO(n11), .S(product[8]) );
  FA_X1 U13 ( .A(a[6]), .B(a[4]), .CI(n13), .CO(n12), .S(product[7]) );
  FA_X1 U14 ( .A(a[5]), .B(a[3]), .CI(n14), .CO(n13), .S(product[6]) );
  FA_X1 U15 ( .A(a[4]), .B(a[2]), .CI(n15), .CO(n14), .S(product[5]) );
  FA_X1 U16 ( .A(a[3]), .B(a[1]), .CI(n16), .CO(n15), .S(product[4]) );
  HA_X1 U17 ( .A(a[0]), .B(a[2]), .CO(n16), .S(product[3]) );
  CLKBUF_X1 U22 ( .A(a[1]), .Z(product[2]) );
  CLKBUF_X1 U23 ( .A(a[0]), .Z(product[1]) );
endmodule


module fir_16tap_DW_mult_uns_2 ( a, b, product );
  input [15:0] a;
  input [3:0] b;
  output [19:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97;

  FA_X1 U6 ( .A(a[12]), .B(n80), .CI(n4), .CO(n3), .S(product[16]) );
  FA_X1 U7 ( .A(a[11]), .B(n81), .CI(n5), .CO(n4), .S(product[15]) );
  FA_X1 U8 ( .A(a[10]), .B(n82), .CI(n6), .CO(n5), .S(product[14]) );
  FA_X1 U9 ( .A(a[9]), .B(n83), .CI(n7), .CO(n6), .S(product[13]) );
  FA_X1 U10 ( .A(a[8]), .B(n84), .CI(n8), .CO(n7), .S(product[12]) );
  FA_X1 U11 ( .A(a[7]), .B(n85), .CI(n9), .CO(n8), .S(product[11]) );
  FA_X1 U12 ( .A(a[6]), .B(n86), .CI(n10), .CO(n9), .S(product[10]) );
  FA_X1 U13 ( .A(a[5]), .B(n87), .CI(n11), .CO(n10), .S(product[9]) );
  FA_X1 U14 ( .A(a[4]), .B(n88), .CI(n12), .CO(n11), .S(product[8]) );
  FA_X1 U15 ( .A(a[3]), .B(n89), .CI(n13), .CO(n12), .S(product[7]) );
  FA_X1 U16 ( .A(a[2]), .B(n90), .CI(n14), .CO(n13), .S(product[6]) );
  FA_X1 U17 ( .A(a[1]), .B(n91), .CI(n15), .CO(n14), .S(product[5]) );
  FA_X1 U18 ( .A(a[0]), .B(n92), .CI(n16), .CO(n15), .S(product[4]) );
  HA_X1 U19 ( .A(n93), .B(n17), .CO(n16), .S(product[3]) );
  HA_X1 U20 ( .A(n94), .B(n95), .CO(n17), .S(product[2]) );
  INV_X1 U42 ( .A(a[1]), .ZN(n94) );
  INV_X1 U43 ( .A(a[0]), .ZN(n95) );
  INV_X1 U44 ( .A(a[2]), .ZN(n93) );
  INV_X1 U45 ( .A(a[3]), .ZN(n92) );
  INV_X1 U46 ( .A(a[15]), .ZN(n80) );
  INV_X1 U47 ( .A(a[4]), .ZN(n91) );
  INV_X1 U48 ( .A(a[5]), .ZN(n90) );
  INV_X1 U49 ( .A(a[6]), .ZN(n89) );
  INV_X1 U50 ( .A(a[7]), .ZN(n88) );
  INV_X1 U51 ( .A(a[8]), .ZN(n87) );
  INV_X1 U52 ( .A(a[9]), .ZN(n86) );
  INV_X1 U53 ( .A(a[10]), .ZN(n85) );
  INV_X1 U54 ( .A(a[11]), .ZN(n84) );
  INV_X1 U55 ( .A(a[12]), .ZN(n83) );
  INV_X1 U56 ( .A(a[13]), .ZN(n82) );
  INV_X1 U57 ( .A(a[14]), .ZN(n81) );
  CLKBUF_X1 U58 ( .A(a[0]), .Z(product[1]) );
  XNOR2_X1 U59 ( .A(a[15]), .B(n96), .ZN(product[19]) );
  NAND2_X1 U60 ( .A1(n97), .A2(n81), .ZN(n96) );
  XNOR2_X1 U61 ( .A(n81), .B(n97), .ZN(product[18]) );
  NOR2_X1 U62 ( .A1(n3), .A2(a[13]), .ZN(n97) );
  XNOR2_X1 U63 ( .A(a[13]), .B(n3), .ZN(product[17]) );
endmodule


module fir_16tap_DW01_add_8 ( A, B, CI, SUM, CO );
  input [21:0] A;
  input [21:0] B;
  output [21:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [19:3] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(SUM[20]), .S(SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n2), .CO(carry[3]), .S(SUM[2]) );
  XOR2_X1 U1 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  AND2_X1 U2 ( .A1(B[1]), .A2(A[1]), .ZN(n2) );
endmodule


module fir_16tap_DW01_add_7 ( A, B, CI, SUM, CO );
  input [22:0] A;
  input [22:0] B;
  output [22:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [20:3] carry;

  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  AND2_X1 U1 ( .A1(B[1]), .A2(A[1]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR2_X1 U3 ( .A(B[20]), .B(carry[20]), .Z(SUM[20]) );
  AND2_X1 U4 ( .A1(B[20]), .A2(carry[20]), .ZN(SUM[21]) );
  CLKBUF_X1 U5 ( .A(A[0]), .Z(SUM[0]) );
endmodule


module fir_16tap_DW01_add_5 ( A, B, CI, SUM, CO );
  input [26:0] A;
  input [26:0] B;
  output [26:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n8;
  wire   [19:3] carry;

  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n2), .CO(carry[3]), .S(SUM[2]) );
  XOR2_X1 U1 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  AND2_X1 U2 ( .A1(B[1]), .A2(A[1]), .ZN(n2) );
  AND2_X1 U3 ( .A1(A[20]), .A2(n8), .ZN(n3) );
  AND2_X1 U4 ( .A1(A[21]), .A2(n3), .ZN(SUM[22]) );
  XOR2_X1 U5 ( .A(A[19]), .B(carry[19]), .Z(SUM[19]) );
  XOR2_X1 U6 ( .A(A[20]), .B(n8), .Z(SUM[20]) );
  XOR2_X1 U7 ( .A(A[21]), .B(n3), .Z(SUM[21]) );
  AND2_X1 U8 ( .A1(A[19]), .A2(carry[19]), .ZN(n8) );
  CLKBUF_X1 U9 ( .A(A[0]), .Z(SUM[0]) );
endmodule


module fir_16tap_DW01_add_4 ( A, B, CI, SUM, CO );
  input [27:0] A;
  input [27:0] B;
  output [27:0] SUM;
  input CI;
  output CO;
  wire   n3;
  wire   [22:2] carry;

  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[22]), .A2(carry[22]), .ZN(SUM[23]) );
  XOR2_X1 U2 ( .A(B[22]), .B(carry[22]), .Z(SUM[22]) );
  AND2_X1 U3 ( .A1(B[0]), .A2(A[0]), .ZN(n3) );
  XOR2_X1 U4 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fir_16tap_DW01_add_3 ( A, B, CI, SUM, CO );
  input [30:0] A;
  input [30:0] B;
  output [30:0] SUM;
  input CI;
  output CO;
  wire   n1, n6;
  wire   [22:2] carry;

  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n6), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[22]), .A2(carry[22]), .ZN(n1) );
  AND2_X1 U2 ( .A1(A[23]), .A2(n1), .ZN(SUM[24]) );
  XOR2_X1 U3 ( .A(A[23]), .B(n1), .Z(SUM[23]) );
  XOR2_X1 U4 ( .A(A[22]), .B(carry[22]), .Z(SUM[22]) );
  XOR2_X1 U5 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U6 ( .A1(B[0]), .A2(A[0]), .ZN(n6) );
endmodule


module fir_16tap_DW_mult_uns_1 ( a, b, product );
  input [15:0] a;
  input [3:0] b;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  HA_X1 U2 ( .A(a[15]), .B(n2), .CO(product[19]), .S(product[18]) );
  FA_X1 U3 ( .A(n19), .B(a[14]), .CI(n3), .CO(n2), .S(product[17]) );
  FA_X1 U4 ( .A(n21), .B(n20), .CI(n4), .CO(n3), .S(product[16]) );
  FA_X1 U5 ( .A(n22), .B(n23), .CI(n5), .CO(n4), .S(product[15]) );
  FA_X1 U6 ( .A(n24), .B(n25), .CI(n6), .CO(n5), .S(product[14]) );
  FA_X1 U7 ( .A(n26), .B(n27), .CI(n7), .CO(n6), .S(product[13]) );
  FA_X1 U8 ( .A(n28), .B(n29), .CI(n8), .CO(n7), .S(product[12]) );
  FA_X1 U9 ( .A(n30), .B(n31), .CI(n9), .CO(n8), .S(product[11]) );
  FA_X1 U10 ( .A(n32), .B(n33), .CI(n10), .CO(n9), .S(product[10]) );
  FA_X1 U11 ( .A(n34), .B(n35), .CI(n11), .CO(n10), .S(product[9]) );
  FA_X1 U12 ( .A(n36), .B(n37), .CI(n12), .CO(n11), .S(product[8]) );
  FA_X1 U13 ( .A(n38), .B(n39), .CI(n13), .CO(n12), .S(product[7]) );
  FA_X1 U14 ( .A(n40), .B(n41), .CI(n14), .CO(n13), .S(product[6]) );
  FA_X1 U15 ( .A(n42), .B(n43), .CI(n15), .CO(n14), .S(product[5]) );
  FA_X1 U16 ( .A(n44), .B(n45), .CI(n16), .CO(n15), .S(product[4]) );
  FA_X1 U17 ( .A(n46), .B(a[0]), .CI(n17), .CO(n16), .S(product[3]) );
  FA_X1 U18 ( .A(a[2]), .B(a[1]), .CI(n18), .CO(n17), .S(product[2]) );
  HA_X1 U19 ( .A(a[0]), .B(a[1]), .CO(n18), .S(product[1]) );
  HA_X1 U20 ( .A(a[15]), .B(a[13]), .CO(n19), .S(n20) );
  FA_X1 U21 ( .A(a[12]), .B(a[15]), .CI(a[14]), .CO(n21), .S(n22) );
  FA_X1 U22 ( .A(a[11]), .B(a[14]), .CI(a[13]), .CO(n23), .S(n24) );
  FA_X1 U23 ( .A(a[10]), .B(a[13]), .CI(a[12]), .CO(n25), .S(n26) );
  FA_X1 U24 ( .A(a[9]), .B(a[12]), .CI(a[11]), .CO(n27), .S(n28) );
  FA_X1 U25 ( .A(a[8]), .B(a[11]), .CI(a[10]), .CO(n29), .S(n30) );
  FA_X1 U26 ( .A(a[7]), .B(a[10]), .CI(a[9]), .CO(n31), .S(n32) );
  FA_X1 U27 ( .A(a[6]), .B(a[9]), .CI(a[8]), .CO(n33), .S(n34) );
  FA_X1 U28 ( .A(a[5]), .B(a[8]), .CI(a[7]), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(a[4]), .B(a[7]), .CI(a[6]), .CO(n37), .S(n38) );
  FA_X1 U30 ( .A(a[3]), .B(a[6]), .CI(a[5]), .CO(n39), .S(n40) );
  FA_X1 U31 ( .A(a[2]), .B(a[5]), .CI(a[4]), .CO(n41), .S(n42) );
  FA_X1 U32 ( .A(a[1]), .B(a[4]), .CI(a[3]), .CO(n43), .S(n44) );
  HA_X1 U33 ( .A(a[3]), .B(a[2]), .CO(n45), .S(n46) );
  CLKBUF_X1 U38 ( .A(a[0]), .Z(product[0]) );
endmodule


module fir_16tap_DW_mult_uns_0 ( a, b, product );
  input [15:0] a;
  input [3:0] b;
  output [19:0] product;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99;

  FA_X1 U8 ( .A(a[11]), .B(n81), .CI(n5), .CO(n4), .S(product[15]) );
  FA_X1 U9 ( .A(a[10]), .B(n82), .CI(n6), .CO(n5), .S(product[14]) );
  FA_X1 U10 ( .A(a[9]), .B(n83), .CI(n7), .CO(n6), .S(product[13]) );
  FA_X1 U11 ( .A(a[8]), .B(n84), .CI(n8), .CO(n7), .S(product[12]) );
  FA_X1 U12 ( .A(a[7]), .B(n85), .CI(n9), .CO(n8), .S(product[11]) );
  FA_X1 U13 ( .A(a[6]), .B(n86), .CI(n10), .CO(n9), .S(product[10]) );
  FA_X1 U14 ( .A(a[5]), .B(n87), .CI(n11), .CO(n10), .S(product[9]) );
  FA_X1 U15 ( .A(a[4]), .B(n88), .CI(n12), .CO(n11), .S(product[8]) );
  FA_X1 U16 ( .A(a[3]), .B(n89), .CI(n13), .CO(n12), .S(product[7]) );
  FA_X1 U17 ( .A(a[2]), .B(n90), .CI(n14), .CO(n13), .S(product[6]) );
  FA_X1 U18 ( .A(a[1]), .B(n91), .CI(n15), .CO(n14), .S(product[5]) );
  FA_X1 U19 ( .A(a[0]), .B(n92), .CI(n16), .CO(n15), .S(product[4]) );
  HA_X1 U20 ( .A(n93), .B(n17), .CO(n16), .S(product[3]) );
  HA_X1 U21 ( .A(n94), .B(n18), .CO(n17), .S(product[2]) );
  HA_X1 U22 ( .A(n95), .B(n96), .CO(n18), .S(product[1]) );
  INV_X1 U43 ( .A(a[1]), .ZN(n95) );
  INV_X1 U44 ( .A(a[0]), .ZN(n96) );
  INV_X1 U45 ( .A(a[2]), .ZN(n94) );
  INV_X1 U46 ( .A(a[3]), .ZN(n93) );
  INV_X1 U47 ( .A(a[4]), .ZN(n92) );
  INV_X1 U48 ( .A(a[5]), .ZN(n91) );
  INV_X1 U49 ( .A(a[6]), .ZN(n90) );
  INV_X1 U50 ( .A(a[7]), .ZN(n89) );
  INV_X1 U51 ( .A(a[8]), .ZN(n88) );
  INV_X1 U52 ( .A(a[9]), .ZN(n87) );
  INV_X1 U53 ( .A(a[10]), .ZN(n86) );
  INV_X1 U54 ( .A(a[11]), .ZN(n85) );
  INV_X1 U55 ( .A(a[12]), .ZN(n84) );
  INV_X1 U56 ( .A(a[13]), .ZN(n83) );
  INV_X1 U57 ( .A(a[15]), .ZN(n81) );
  INV_X1 U58 ( .A(a[14]), .ZN(n82) );
  CLKBUF_X1 U59 ( .A(a[0]), .Z(product[0]) );
  XOR2_X1 U60 ( .A(n81), .B(n97), .Z(product[19]) );
  NAND2_X1 U61 ( .A1(n98), .A2(n82), .ZN(n97) );
  XOR2_X1 U62 ( .A(a[14]), .B(n98), .Z(product[18]) );
  NOR2_X1 U63 ( .A1(n99), .A2(a[13]), .ZN(n98) );
  XOR2_X1 U64 ( .A(n83), .B(n99), .Z(product[17]) );
  OR2_X1 U65 ( .A1(n4), .A2(a[12]), .ZN(n99) );
  XOR2_X1 U66 ( .A(n84), .B(n4), .Z(product[16]) );
endmodule


module fir_16tap_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n7, n9;
  wire   [21:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n9), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[22]), .A2(n7), .ZN(n1) );
  AND2_X1 U2 ( .A1(B[23]), .A2(n1), .ZN(n2) );
  AND2_X1 U3 ( .A1(B[24]), .A2(n2), .ZN(SUM[25]) );
  XOR2_X1 U4 ( .A(B[22]), .B(n7), .Z(SUM[22]) );
  XOR2_X1 U5 ( .A(B[23]), .B(n1), .Z(SUM[23]) );
  XOR2_X1 U6 ( .A(B[24]), .B(n2), .Z(SUM[24]) );
  AND2_X1 U7 ( .A1(B[21]), .A2(carry[21]), .ZN(n7) );
  XOR2_X1 U8 ( .A(B[21]), .B(carry[21]), .Z(SUM[21]) );
  AND2_X1 U9 ( .A1(B[0]), .A2(A[0]), .ZN(n9) );
  XOR2_X1 U10 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fir_16tap_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n9, n11, n12, n15, n16, n19, n21;
  wire   [16:2] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n21), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(A[22]), .A2(n9), .ZN(n1) );
  AND2_X1 U2 ( .A1(A[23]), .A2(n1), .ZN(n2) );
  AND2_X1 U3 ( .A1(A[24]), .A2(n2), .ZN(n3) );
  XOR2_X1 U4 ( .A(A[25]), .B(n3), .Z(SUM[25]) );
  XOR2_X1 U5 ( .A(A[22]), .B(n9), .Z(SUM[22]) );
  XOR2_X1 U6 ( .A(A[23]), .B(n1), .Z(SUM[23]) );
  XOR2_X1 U7 ( .A(A[24]), .B(n2), .Z(SUM[24]) );
  AND2_X1 U8 ( .A1(A[25]), .A2(n3), .ZN(SUM[26]) );
  AND2_X1 U9 ( .A1(A[21]), .A2(n12), .ZN(n9) );
  XOR2_X1 U10 ( .A(A[21]), .B(n12), .Z(SUM[21]) );
  AND2_X1 U11 ( .A1(A[19]), .A2(n16), .ZN(n11) );
  AND2_X1 U12 ( .A1(A[20]), .A2(n11), .ZN(n12) );
  XOR2_X1 U13 ( .A(A[19]), .B(n16), .Z(SUM[19]) );
  XOR2_X1 U14 ( .A(A[20]), .B(n11), .Z(SUM[20]) );
  AND2_X1 U15 ( .A1(A[17]), .A2(n19), .ZN(n15) );
  AND2_X1 U16 ( .A1(A[18]), .A2(n15), .ZN(n16) );
  XOR2_X1 U17 ( .A(A[18]), .B(n15), .Z(SUM[18]) );
  XOR2_X1 U18 ( .A(A[17]), .B(n19), .Z(SUM[17]) );
  AND2_X1 U19 ( .A1(A[16]), .A2(carry[16]), .ZN(n19) );
  XOR2_X1 U20 ( .A(A[16]), .B(carry[16]), .Z(SUM[16]) );
  AND2_X1 U21 ( .A1(B[0]), .A2(A[0]), .ZN(n21) );
  XOR2_X1 U22 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fir_16tap ( x, clk, reset, y );
  input [15:0] x;
  output [31:0] y;
  input clk, reset;
  wire   m43_9_, m43_8_, m43_7_, m43_6_, m43_5_, m43_4_, m43_3_, m43_2_,
         m43_20_, m43_1_, m43_19_, m43_18_, m43_17_, m43_16_, m43_15_, m43_14_,
         m43_13_, m43_12_, m43_11_, m43_10_, m43_0_, m42_9_, m42_8_, m42_7_,
         m42_6_, m42_5_, m42_4_, m42_3_, m42_2_, m42_1_, m42_19_, m42_18_,
         m42_17_, m42_16_, m42_15_, m42_14_, m42_13_, m42_12_, m42_11_,
         m42_10_, m42_0_, m40_9_, m40_8_, m40_7_, m40_6_, m40_5_, m40_4_,
         m40_3_, m40_2_, m40_1_, m40_19_, m40_18_, m40_17_, m40_16_, m40_15_,
         m40_14_, m40_13_, m40_12_, m40_11_, m40_10_, m39_9_, m39_8_, m39_7_,
         m39_6_, m39_5_, m39_4_, m39_3_, m39_2_, m39_1_, m39_19_, m39_18_,
         m39_17_, m39_16_, m39_15_, m39_14_, m39_13_, m39_12_, m39_11_,
         m39_10_, m39_0_, m38_9_, m38_8_, m38_7_, m38_6_, m38_5_, m38_4_,
         m38_3_, m38_2_, m38_1_, m38_19_, m38_18_, m38_17_, m38_16_, m38_15_,
         m38_14_, m38_13_, m38_12_, m38_11_, m38_10_, m38_0_, m37_9_, m37_8_,
         m37_7_, m37_6_, m37_5_, m37_4_, m37_3_, m37_2_, m37_20_, m37_1_,
         m37_19_, m37_18_, m37_17_, m37_16_, m37_15_, m37_14_, m37_13_,
         m37_12_, m37_11_, m37_10_, m37_0_, m36_9_, m36_8_, m36_7_, m36_6_,
         m36_5_, m36_4_, m36_3_, m36_2_, m36_19_, m36_18_, m36_17_, m36_16_,
         m36_15_, m36_14_, m36_13_, m36_12_, m36_11_, m36_10_, m35_9_, m35_8_,
         m35_7_, m35_6_, m35_5_, m35_4_, m35_3_, m35_2_, m35_22_, m35_21_,
         m35_20_, m35_1_, m35_19_, m35_18_, m35_17_, m35_16_, m35_15_, m35_14_,
         m35_13_, m35_12_, m35_11_, m35_10_, m35_0_, m34_9_, m34_8_, m34_7_,
         m34_6_, m34_5_, m34_4_, m34_3_, m34_2_, m34_1_, m34_19_, m34_18_,
         m34_17_, m34_16_, m34_15_, m34_14_, m34_13_, m34_12_, m34_11_,
         m34_10_, m34_0_, m32_9_, m32_8_, m32_7_, m32_6_, m32_5_, m32_4_,
         m32_3_, m32_2_, m32_1_, m32_19_, m32_18_, m32_17_, m32_16_, m32_15_,
         m32_14_, m32_13_, m32_12_, m32_11_, m32_10_, m31_9_, m31_8_, m31_7_,
         m31_6_, m31_5_, m31_4_, m31_3_, m31_2_, m31_1_, m31_18_, m31_17_,
         m31_16_, m31_15_, m31_14_, m31_13_, m31_12_, m31_11_, m31_10_, m30_9_,
         m30_8_, m30_7_, m30_6_, m30_5_, m30_4_, m30_3_, m30_2_, m30_19_,
         m30_18_, m30_17_, m30_16_, m30_15_, m30_14_, m30_13_, m30_12_,
         m30_11_, m30_10_, m29_9_, m29_8_, m29_7_, m29_6_, m29_5_, m29_4_,
         m29_3_, m29_20_, m29_19_, m29_18_, m29_17_, m29_16_, m29_15_, m29_14_,
         m29_13_, m29_12_, m29_11_, m29_10_, m27_9_, m27_8_, m27_7_, m27_6_,
         m27_5_, m27_4_, m27_3_, m27_2_, m27_1_, m27_19_, m27_18_, m27_17_,
         m27_16_, m27_15_, m27_14_, m27_13_, m27_12_, m27_11_, m27_10_, m27_0_,
         m26_9_, m26_8_, m26_7_, m26_6_, m26_5_, m26_4_, m26_3_, m26_2_,
         m26_1_, m26_18_, m26_17_, m26_16_, m26_15_, m26_14_, m26_13_, m26_12_,
         m26_11_, m26_10_, m26_0_, m25_9_, m25_8_, m25_7_, m25_6_, m25_5_,
         m25_4_, m25_3_, m25_2_, m25_20_, m25_1_, m25_19_, m25_18_, m25_17_,
         m25_16_, m25_15_, m25_14_, m25_13_, m25_12_, m25_11_, m25_10_, m24_9_,
         m24_8_, m24_7_, m24_6_, m24_5_, m24_4_, m24_3_, m24_2_, m24_1_,
         m24_18_, m24_17_, m24_16_, m24_15_, m24_14_, m24_13_, m24_12_,
         m24_11_, m24_10_, m22_9_, m22_8_, m22_7_, m22_6_, m22_5_, m22_4_,
         m22_3_, m22_2_, m22_1_, m22_18_, m22_17_, m22_16_, m22_15_, m22_14_,
         m22_13_, m22_12_, m22_11_, m22_10_, m22_0_, m18_9_, m18_8_, m18_7_,
         m18_6_, m18_5_, m18_4_, m18_3_, m18_2_, m18_1_, m18_17_, m18_16_,
         m18_15_, m18_14_, m18_13_, m18_12_, m18_11_, m18_10_,
         add_6_root_add_0_root_add_94_carry_4_,
         add_6_root_add_0_root_add_94_carry_5_,
         add_6_root_add_0_root_add_94_carry_6_,
         add_6_root_add_0_root_add_94_carry_7_,
         add_6_root_add_0_root_add_94_carry_8_,
         add_6_root_add_0_root_add_94_carry_9_,
         add_6_root_add_0_root_add_94_carry_10_,
         add_6_root_add_0_root_add_94_carry_11_,
         add_6_root_add_0_root_add_94_carry_12_,
         add_6_root_add_0_root_add_94_carry_13_,
         add_6_root_add_0_root_add_94_carry_14_,
         add_6_root_add_0_root_add_94_carry_15_,
         add_6_root_add_0_root_add_94_carry_16_,
         add_6_root_add_0_root_add_94_carry_17_,
         add_6_root_add_0_root_add_94_carry_18_,
         add_6_root_add_0_root_add_94_carry_19_,
         add_6_root_add_0_root_add_94_carry_20_,
         add_6_root_add_0_root_add_94_carry_21_,
         add_6_root_add_0_root_add_94_SUM_3_,
         add_6_root_add_0_root_add_94_SUM_4_,
         add_6_root_add_0_root_add_94_SUM_5_,
         add_6_root_add_0_root_add_94_SUM_6_,
         add_6_root_add_0_root_add_94_SUM_7_,
         add_6_root_add_0_root_add_94_SUM_8_,
         add_6_root_add_0_root_add_94_SUM_9_,
         add_6_root_add_0_root_add_94_SUM_10_,
         add_6_root_add_0_root_add_94_SUM_11_,
         add_6_root_add_0_root_add_94_SUM_12_,
         add_6_root_add_0_root_add_94_SUM_13_,
         add_6_root_add_0_root_add_94_SUM_14_,
         add_6_root_add_0_root_add_94_SUM_15_,
         add_6_root_add_0_root_add_94_SUM_16_,
         add_6_root_add_0_root_add_94_SUM_17_,
         add_6_root_add_0_root_add_94_SUM_18_,
         add_6_root_add_0_root_add_94_SUM_19_,
         add_6_root_add_0_root_add_94_SUM_20_, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44;
  wire   [15:1] m0;
  wire   [15:0] m1;
  wire   [15:0] m2;
  wire   [15:0] m3;
  wire   [15:0] m4;
  wire   [15:0] m5;
  wire   [15:1] m6;
  wire   [15:0] m7;
  wire   [15:0] m8;
  wire   [15:0] m9;
  wire   [15:0] m10;
  wire   [15:0] m11;
  wire   [15:0] m12;
  wire   [15:0] m13;
  wire   [15:0] m14;
  wire   [19:1] add_8_root_add_0_root_add_94_carry;
  wire   [17:3] add_14_root_add_0_root_add_94_carry;
  wire   [19:5] add_13_root_add_0_root_add_94_carry;
  wire   [18:2] add_12_root_add_0_root_add_94_carry;
  wire   [19:3] add_9_root_add_0_root_add_94_carry;

  dff_16bit_0 q1 ( .d(x), .clk(clk), .reset(reset), .q({m0, m31_1_}) );
  dff_16bit_14 q2 ( .d({m0, m31_1_}), .clk(clk), .reset(reset), .q(m1) );
  dff_16bit_13 q3 ( .d(m1), .clk(clk), .reset(reset), .q(m2) );
  dff_16bit_12 q4 ( .d(m2), .clk(clk), .reset(reset), .q(m3) );
  dff_16bit_11 q5 ( .d(m3), .clk(clk), .reset(reset), .q(m4) );
  dff_16bit_10 q6 ( .d(m4), .clk(clk), .reset(reset), .q(m5) );
  dff_16bit_9 q7 ( .d(m5), .clk(clk), .reset(reset), .q({m6, m29_3_}) );
  dff_16bit_8 q8 ( .d({m6, m29_3_}), .clk(clk), .reset(reset), .q(m7) );
  dff_16bit_7 q9 ( .d(m7), .clk(clk), .reset(reset), .q(m8) );
  dff_16bit_6 q10 ( .d(m8), .clk(clk), .reset(reset), .q(m9) );
  dff_16bit_5 q11 ( .d(m9), .clk(clk), .reset(reset), .q(m10) );
  dff_16bit_4 q12 ( .d(m10), .clk(clk), .reset(reset), .q(m11) );
  dff_16bit_3 q13 ( .d(m11), .clk(clk), .reset(reset), .q(m12) );
  dff_16bit_2 q14 ( .d(m12), .clk(clk), .reset(reset), .q(m13) );
  dff_16bit_1 q15 ( .d(m13), .clk(clk), .reset(reset), .q(m14) );
  fir_16tap_DW_mult_uns_10 mult_73 ( .a(m10), .b({1'b1, 1'b1, 1'b0, 1'b0}), 
        .product({m36_19_, m36_18_, m36_17_, m36_16_, m36_15_, m36_14_, 
        m36_13_, m36_12_, m36_11_, m36_10_, m36_9_, m36_8_, m36_7_, m36_6_, 
        m36_5_, m36_4_, m36_3_, m36_2_, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}) );
  fir_16tap_DW_mult_uns_9 mult_70 ( .a(m7), .b({1'b1, 1'b0, 1'b0, 1'b1}), 
        .product({m30_19_, m30_18_, m30_17_, m30_16_, m30_15_, m30_14_, 
        m30_13_, m30_12_, m30_11_, m30_10_, m30_9_, m30_8_, m30_7_, m30_6_, 
        m30_5_, m30_4_, m30_3_, m30_2_, m37_1_, m37_0_}) );
  fir_16tap_DW_mult_uns_8 mult_64 ( .a(m1), .b({1'b1, 1'b1}), .product({
        m18_17_, m18_16_, m18_15_, m18_14_, m18_13_, m18_12_, m18_11_, m18_10_, 
        m18_9_, m18_8_, m18_7_, m18_6_, m18_5_, m18_4_, m18_3_, m18_2_, m18_1_, 
        m39_0_}) );
  fir_16tap_DW_mult_uns_7 mult_67 ( .a(m4), .b({1'b1, 1'b1, 1'b0}), .product({
        m24_18_, m24_17_, m24_16_, m24_15_, m24_14_, m24_13_, m24_12_, m24_11_, 
        m24_10_, m24_9_, m24_8_, m24_7_, m24_6_, m24_5_, m24_4_, m24_3_, 
        m24_2_, m24_1_, SYNOPSYS_UNCONNECTED_3}) );
  fir_16tap_DW01_add_12 add_3_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m37_20_, m37_19_, m37_18_, m37_17_, 
        m37_16_, m37_15_, m37_14_, m37_13_, m37_12_, m37_11_, m37_10_, m37_9_, 
        m37_8_, m37_7_, m37_6_, m37_5_, m37_4_, m37_3_, m37_2_, m37_1_, m37_0_}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m39_19_, 
        m39_18_, m39_17_, m39_16_, m39_15_, m39_14_, m39_13_, m39_12_, m39_11_, 
        m39_10_, m39_9_, m39_8_, m39_7_, m39_6_, m39_5_, m39_4_, m39_3_, 
        m39_2_, m39_1_, m39_0_}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69, n68, n67, n66, n65, n64, 
        n63, n62, n61, n60}) );
  fir_16tap_DW_mult_uns_6 mult_68 ( .a(m5), .b({1'b1, 1'b1, 1'b1}), .product({
        m26_18_, m26_17_, m26_16_, m26_15_, m26_14_, m26_13_, m26_12_, m26_11_, 
        m26_10_, m26_9_, m26_8_, m26_7_, m26_6_, m26_5_, m26_4_, m26_3_, 
        m26_2_, m26_1_, m26_0_}) );
  fir_16tap_DW_mult_uns_5 mult_66 ( .a(m3), .b({1'b1, 1'b0, 1'b1}), .product({
        m22_18_, m22_17_, m22_16_, m22_15_, m22_14_, m22_13_, m22_12_, m22_11_, 
        m22_10_, m22_9_, m22_8_, m22_7_, m22_6_, m22_5_, m22_4_, m22_3_, 
        m22_2_, m22_1_, m22_0_}) );
  fir_16tap_DW01_add_11 add_11_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, m26_18_, m26_17_, m26_16_, m26_15_, m26_14_, m26_13_, m26_12_, 
        m26_11_, m26_10_, m26_9_, m26_8_, m26_7_, m26_6_, m26_5_, m26_4_, 
        m26_3_, m26_2_, m26_1_, m26_0_}), .B({1'b0, 1'b0, 1'b0, 1'b0, m22_18_, 
        m22_17_, m22_16_, m22_15_, m22_14_, m22_13_, m22_12_, m22_11_, m22_10_, 
        m22_9_, m22_8_, m22_7_, m22_6_, m22_5_, m22_4_, m22_3_, m22_2_, m22_1_, 
        m22_0_}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, m27_19_, m27_18_, 
        m27_17_, m27_16_, m27_15_, m27_14_, m27_13_, m27_12_, m27_11_, m27_10_, 
        m27_9_, m27_8_, m27_7_, m27_6_, m27_5_, m27_4_, m27_3_, m27_2_, m27_1_, 
        m27_0_}) );
  fir_16tap_DW_mult_uns_4 mult_74 ( .a(m11), .b({1'b1, 1'b1, 1'b0, 1'b1}), 
        .product({m38_19_, m38_18_, m38_17_, m38_16_, m38_15_, m38_14_, 
        m38_13_, m38_12_, m38_11_, m38_10_, m38_9_, m38_8_, m38_7_, m38_6_, 
        m38_5_, m38_4_, m38_3_, m38_2_, m38_1_, m38_0_}) );
  fir_16tap_DW_mult_uns_3 mult_71 ( .a(m8), .b({1'b1, 1'b0, 1'b1, 1'b0}), 
        .product({m32_19_, m32_18_, m32_17_, m32_16_, m32_15_, m32_14_, 
        m32_13_, m32_12_, m32_11_, m32_10_, m32_9_, m32_8_, m32_7_, m32_6_, 
        m32_5_, m32_4_, m32_3_, m32_2_, m32_1_, SYNOPSYS_UNCONNECTED_15}) );
  fir_16tap_DW_mult_uns_2 mult_75 ( .a(m12), .b({1'b1, 1'b1, 1'b1, 1'b0}), 
        .product({m40_19_, m40_18_, m40_17_, m40_16_, m40_15_, m40_14_, 
        m40_13_, m40_12_, m40_11_, m40_10_, m40_9_, m40_8_, m40_7_, m40_6_, 
        m40_5_, m40_4_, m40_3_, m40_2_, m40_1_, SYNOPSYS_UNCONNECTED_16}) );
  fir_16tap_DW01_add_8 add_10_root_add_0_root_add_94 ( .A({1'b0, 1'b0, m32_19_, 
        m32_18_, m32_17_, m32_16_, m32_15_, m32_14_, m32_13_, m32_12_, m32_11_, 
        m32_10_, m32_9_, m32_8_, m32_7_, m32_6_, m32_5_, m32_4_, m32_3_, 
        m32_2_, m32_1_, 1'b0}), .B({1'b0, 1'b0, m40_19_, m40_18_, m40_17_, 
        m40_16_, m40_15_, m40_14_, m40_13_, m40_12_, m40_11_, m40_10_, m40_9_, 
        m40_8_, m40_7_, m40_6_, m40_5_, m40_4_, m40_3_, m40_2_, m40_1_, 1'b0}), 
        .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED_17, m25_20_, m25_19_, m25_18_, 
        m25_17_, m25_16_, m25_15_, m25_14_, m25_13_, m25_12_, m25_11_, m25_10_, 
        m25_9_, m25_8_, m25_7_, m25_6_, m25_5_, m25_4_, m25_3_, m25_2_, m25_1_, 
        SYNOPSYS_UNCONNECTED_18}) );
  fir_16tap_DW01_add_7 add_7_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        m38_19_, m38_18_, m38_17_, m38_16_, m38_15_, m38_14_, m38_13_, m38_12_, 
        m38_11_, m38_10_, m38_9_, m38_8_, m38_7_, m38_6_, m38_5_, m38_4_, 
        m38_3_, m38_2_, m38_1_, m38_0_}), .B({1'b0, 1'b0, m25_20_, m25_19_, 
        m25_18_, m25_17_, m25_16_, m25_15_, m25_14_, m25_13_, m25_12_, m25_11_, 
        m25_10_, m25_9_, m25_8_, m25_7_, m25_6_, m25_5_, m25_4_, m25_3_, 
        m25_2_, m25_1_, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED_19, n35, 
        n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, n21, 
        n20, n19, n18, n17, n16, n15, n14}) );
  fir_16tap_DW01_add_5 add_5_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, n35, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, 
        n23, n22, n21, n20, n19, n18, n17, n16, n15, n14}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m31_18_, m31_17_, m31_16_, m31_15_, 
        m31_14_, m31_13_, m31_12_, m31_11_, m31_10_, m31_9_, m31_8_, m31_7_, 
        m31_6_, m31_5_, m31_4_, m31_3_, m31_2_, m31_1_, 1'b0}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, m35_22_, m35_21_, 
        m35_20_, m35_19_, m35_18_, m35_17_, m35_16_, m35_15_, m35_14_, m35_13_, 
        m35_12_, m35_11_, m35_10_, m35_9_, m35_8_, m35_7_, m35_6_, m35_5_, 
        m35_4_, m35_3_, m35_2_, m35_1_, m35_0_}) );
  fir_16tap_DW01_add_4 add_4_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, add_6_root_add_0_root_add_94_carry_21_, 
        add_6_root_add_0_root_add_94_SUM_20_, 
        add_6_root_add_0_root_add_94_SUM_19_, 
        add_6_root_add_0_root_add_94_SUM_18_, 
        add_6_root_add_0_root_add_94_SUM_17_, 
        add_6_root_add_0_root_add_94_SUM_16_, 
        add_6_root_add_0_root_add_94_SUM_15_, 
        add_6_root_add_0_root_add_94_SUM_14_, 
        add_6_root_add_0_root_add_94_SUM_13_, 
        add_6_root_add_0_root_add_94_SUM_12_, 
        add_6_root_add_0_root_add_94_SUM_11_, 
        add_6_root_add_0_root_add_94_SUM_10_, 
        add_6_root_add_0_root_add_94_SUM_9_, 
        add_6_root_add_0_root_add_94_SUM_8_, 
        add_6_root_add_0_root_add_94_SUM_7_, 
        add_6_root_add_0_root_add_94_SUM_6_, 
        add_6_root_add_0_root_add_94_SUM_5_, 
        add_6_root_add_0_root_add_94_SUM_4_, 
        add_6_root_add_0_root_add_94_SUM_3_, m27_2_, m27_1_, m27_0_}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m35_22_, m35_21_, m35_20_, m35_19_, 
        m35_18_, m35_17_, m35_16_, m35_15_, m35_14_, m35_13_, m35_12_, m35_11_, 
        m35_10_, m35_9_, m35_8_, m35_7_, m35_6_, m35_5_, m35_4_, m35_3_, 
        m35_2_, m35_1_, m35_0_}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, n59, n58, n57, n56, n55, n54, n53, n52, n51, 
        n50, n49, n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, 
        n36}) );
  fir_16tap_DW01_add_3 add_2_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, n59, n58, n57, n56, n55, n54, n53, n52, n51, 
        n50, n49, n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, 
        n36}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n81, 
        n80, n79, n78, n77, n76, n75, n74, n73, n72, n71, n70, n69, n68, n67, 
        n66, n65, n64, n63, n62, n61, n60}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, n106, n105, n104, 
        n103, n102, n101, n100, n99, n98, n97, n96, n95, n94, n93, n92, n91, 
        n90, n89, n88, n87, n86, n85, n84, n83, n82}) );
  fir_16tap_DW_mult_uns_1 mult_72 ( .a(m9), .b({1'b1, 1'b0, 1'b1, 1'b1}), 
        .product({m34_19_, m34_18_, m34_17_, m34_16_, m34_15_, m34_14_, 
        m34_13_, m34_12_, m34_11_, m34_10_, m34_9_, m34_8_, m34_7_, m34_6_, 
        m34_5_, m34_4_, m34_3_, m34_2_, m34_1_, m34_0_}) );
  fir_16tap_DW_mult_uns_0 mult_76 ( .a(m13), .b({1'b1, 1'b1, 1'b1, 1'b1}), 
        .product({m42_19_, m42_18_, m42_17_, m42_16_, m42_15_, m42_14_, 
        m42_13_, m42_12_, m42_11_, m42_10_, m42_9_, m42_8_, m42_7_, m42_6_, 
        m42_5_, m42_4_, m42_3_, m42_2_, m42_1_, m42_0_}) );
  fir_16tap_DW01_add_1 add_1_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, m43_20_, m43_19_, 
        m43_18_, m43_17_, m43_16_, m43_15_, m43_14_, m43_13_, m43_12_, m43_11_, 
        m43_10_, m43_9_, m43_8_, m43_7_, m43_6_, m43_5_, m43_4_, m43_3_, 
        m43_2_, m43_1_, m43_0_}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n106, n105, n104, n103, n102, n101, n100, n99, n98, n97, n96, n95, n94, 
        n93, n92, n91, n90, n89, n88, n87, n86, n85, n84, n83, n82}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, n132, n131, n130, 
        n129, n128, n127, n126, n125, n124, n123, n122, n121, n120, n119, n118, 
        n117, n116, n115, n114, n113, n112, n111, n110, n109, n108, n107}) );
  fir_16tap_DW01_add_0 add_0_root_add_0_root_add_94 ( .A({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n132, n131, n130, n129, n128, n127, n126, n125, n124, 
        n123, n122, n121, n120, n119, n118, n117, n116, n115, n114, n113, n112, 
        n111, n110, n109, n108, n107}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, x}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, y[26:0]}) );
  FA_X1 add_8_root_add_0_root_add_94_U1_1 ( .A(m34_1_), .B(m42_1_), .CI(
        add_8_root_add_0_root_add_94_carry[1]), .CO(
        add_8_root_add_0_root_add_94_carry[2]), .S(m43_1_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_2 ( .A(m34_2_), .B(m42_2_), .CI(
        add_8_root_add_0_root_add_94_carry[2]), .CO(
        add_8_root_add_0_root_add_94_carry[3]), .S(m43_2_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_3 ( .A(m34_3_), .B(m42_3_), .CI(
        add_8_root_add_0_root_add_94_carry[3]), .CO(
        add_8_root_add_0_root_add_94_carry[4]), .S(m43_3_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_4 ( .A(m34_4_), .B(m42_4_), .CI(
        add_8_root_add_0_root_add_94_carry[4]), .CO(
        add_8_root_add_0_root_add_94_carry[5]), .S(m43_4_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_5 ( .A(m34_5_), .B(m42_5_), .CI(
        add_8_root_add_0_root_add_94_carry[5]), .CO(
        add_8_root_add_0_root_add_94_carry[6]), .S(m43_5_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_6 ( .A(m34_6_), .B(m42_6_), .CI(
        add_8_root_add_0_root_add_94_carry[6]), .CO(
        add_8_root_add_0_root_add_94_carry[7]), .S(m43_6_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_7 ( .A(m34_7_), .B(m42_7_), .CI(
        add_8_root_add_0_root_add_94_carry[7]), .CO(
        add_8_root_add_0_root_add_94_carry[8]), .S(m43_7_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_8 ( .A(m34_8_), .B(m42_8_), .CI(
        add_8_root_add_0_root_add_94_carry[8]), .CO(
        add_8_root_add_0_root_add_94_carry[9]), .S(m43_8_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_9 ( .A(m34_9_), .B(m42_9_), .CI(
        add_8_root_add_0_root_add_94_carry[9]), .CO(
        add_8_root_add_0_root_add_94_carry[10]), .S(m43_9_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_10 ( .A(m34_10_), .B(m42_10_), .CI(
        add_8_root_add_0_root_add_94_carry[10]), .CO(
        add_8_root_add_0_root_add_94_carry[11]), .S(m43_10_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_11 ( .A(m34_11_), .B(m42_11_), .CI(
        add_8_root_add_0_root_add_94_carry[11]), .CO(
        add_8_root_add_0_root_add_94_carry[12]), .S(m43_11_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_12 ( .A(m34_12_), .B(m42_12_), .CI(
        add_8_root_add_0_root_add_94_carry[12]), .CO(
        add_8_root_add_0_root_add_94_carry[13]), .S(m43_12_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_13 ( .A(m34_13_), .B(m42_13_), .CI(
        add_8_root_add_0_root_add_94_carry[13]), .CO(
        add_8_root_add_0_root_add_94_carry[14]), .S(m43_13_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_14 ( .A(m34_14_), .B(m42_14_), .CI(
        add_8_root_add_0_root_add_94_carry[14]), .CO(
        add_8_root_add_0_root_add_94_carry[15]), .S(m43_14_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_15 ( .A(m34_15_), .B(m42_15_), .CI(
        add_8_root_add_0_root_add_94_carry[15]), .CO(
        add_8_root_add_0_root_add_94_carry[16]), .S(m43_15_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_16 ( .A(m34_16_), .B(m42_16_), .CI(
        add_8_root_add_0_root_add_94_carry[16]), .CO(
        add_8_root_add_0_root_add_94_carry[17]), .S(m43_16_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_17 ( .A(m34_17_), .B(m42_17_), .CI(
        add_8_root_add_0_root_add_94_carry[17]), .CO(
        add_8_root_add_0_root_add_94_carry[18]), .S(m43_17_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_18 ( .A(m34_18_), .B(m42_18_), .CI(
        add_8_root_add_0_root_add_94_carry[18]), .CO(
        add_8_root_add_0_root_add_94_carry[19]), .S(m43_18_) );
  FA_X1 add_8_root_add_0_root_add_94_U1_19 ( .A(m34_19_), .B(m42_19_), .CI(
        add_8_root_add_0_root_add_94_carry[19]), .CO(m43_20_), .S(m43_19_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_3 ( .A(m0[2]), .B(m2[1]), .CI(
        add_14_root_add_0_root_add_94_carry[3]), .CO(
        add_14_root_add_0_root_add_94_carry[4]), .S(m31_3_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_4 ( .A(m0[3]), .B(m2[2]), .CI(
        add_14_root_add_0_root_add_94_carry[4]), .CO(
        add_14_root_add_0_root_add_94_carry[5]), .S(m31_4_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_5 ( .A(m0[4]), .B(m2[3]), .CI(
        add_14_root_add_0_root_add_94_carry[5]), .CO(
        add_14_root_add_0_root_add_94_carry[6]), .S(m31_5_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_6 ( .A(m0[5]), .B(m2[4]), .CI(
        add_14_root_add_0_root_add_94_carry[6]), .CO(
        add_14_root_add_0_root_add_94_carry[7]), .S(m31_6_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_7 ( .A(m0[6]), .B(m2[5]), .CI(
        add_14_root_add_0_root_add_94_carry[7]), .CO(
        add_14_root_add_0_root_add_94_carry[8]), .S(m31_7_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_8 ( .A(m0[7]), .B(m2[6]), .CI(
        add_14_root_add_0_root_add_94_carry[8]), .CO(
        add_14_root_add_0_root_add_94_carry[9]), .S(m31_8_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_9 ( .A(m0[8]), .B(m2[7]), .CI(
        add_14_root_add_0_root_add_94_carry[9]), .CO(
        add_14_root_add_0_root_add_94_carry[10]), .S(m31_9_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_10 ( .A(m0[9]), .B(m2[8]), .CI(
        add_14_root_add_0_root_add_94_carry[10]), .CO(
        add_14_root_add_0_root_add_94_carry[11]), .S(m31_10_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_11 ( .A(m0[10]), .B(m2[9]), .CI(
        add_14_root_add_0_root_add_94_carry[11]), .CO(
        add_14_root_add_0_root_add_94_carry[12]), .S(m31_11_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_12 ( .A(m0[11]), .B(m2[10]), .CI(
        add_14_root_add_0_root_add_94_carry[12]), .CO(
        add_14_root_add_0_root_add_94_carry[13]), .S(m31_12_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_13 ( .A(m0[12]), .B(m2[11]), .CI(
        add_14_root_add_0_root_add_94_carry[13]), .CO(
        add_14_root_add_0_root_add_94_carry[14]), .S(m31_13_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_14 ( .A(m0[13]), .B(m2[12]), .CI(
        add_14_root_add_0_root_add_94_carry[14]), .CO(
        add_14_root_add_0_root_add_94_carry[15]), .S(m31_14_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_15 ( .A(m0[14]), .B(m2[13]), .CI(
        add_14_root_add_0_root_add_94_carry[15]), .CO(
        add_14_root_add_0_root_add_94_carry[16]), .S(m31_15_) );
  FA_X1 add_14_root_add_0_root_add_94_U1_16 ( .A(m0[15]), .B(m2[14]), .CI(
        add_14_root_add_0_root_add_94_carry[16]), .CO(
        add_14_root_add_0_root_add_94_carry[17]), .S(m31_16_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_4 ( .A(m27_4_), .B(m29_4_), .CI(
        add_6_root_add_0_root_add_94_carry_4_), .CO(
        add_6_root_add_0_root_add_94_carry_5_), .S(
        add_6_root_add_0_root_add_94_SUM_4_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_5 ( .A(m27_5_), .B(m29_5_), .CI(
        add_6_root_add_0_root_add_94_carry_5_), .CO(
        add_6_root_add_0_root_add_94_carry_6_), .S(
        add_6_root_add_0_root_add_94_SUM_5_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_6 ( .A(m27_6_), .B(m29_6_), .CI(
        add_6_root_add_0_root_add_94_carry_6_), .CO(
        add_6_root_add_0_root_add_94_carry_7_), .S(
        add_6_root_add_0_root_add_94_SUM_6_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_7 ( .A(m27_7_), .B(m29_7_), .CI(
        add_6_root_add_0_root_add_94_carry_7_), .CO(
        add_6_root_add_0_root_add_94_carry_8_), .S(
        add_6_root_add_0_root_add_94_SUM_7_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_8 ( .A(m27_8_), .B(m29_8_), .CI(
        add_6_root_add_0_root_add_94_carry_8_), .CO(
        add_6_root_add_0_root_add_94_carry_9_), .S(
        add_6_root_add_0_root_add_94_SUM_8_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_9 ( .A(m27_9_), .B(m29_9_), .CI(
        add_6_root_add_0_root_add_94_carry_9_), .CO(
        add_6_root_add_0_root_add_94_carry_10_), .S(
        add_6_root_add_0_root_add_94_SUM_9_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_10 ( .A(m27_10_), .B(m29_10_), .CI(
        add_6_root_add_0_root_add_94_carry_10_), .CO(
        add_6_root_add_0_root_add_94_carry_11_), .S(
        add_6_root_add_0_root_add_94_SUM_10_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_11 ( .A(m27_11_), .B(m29_11_), .CI(
        add_6_root_add_0_root_add_94_carry_11_), .CO(
        add_6_root_add_0_root_add_94_carry_12_), .S(
        add_6_root_add_0_root_add_94_SUM_11_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_12 ( .A(m27_12_), .B(m29_12_), .CI(
        add_6_root_add_0_root_add_94_carry_12_), .CO(
        add_6_root_add_0_root_add_94_carry_13_), .S(
        add_6_root_add_0_root_add_94_SUM_12_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_13 ( .A(m27_13_), .B(m29_13_), .CI(
        add_6_root_add_0_root_add_94_carry_13_), .CO(
        add_6_root_add_0_root_add_94_carry_14_), .S(
        add_6_root_add_0_root_add_94_SUM_13_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_14 ( .A(m27_14_), .B(m29_14_), .CI(
        add_6_root_add_0_root_add_94_carry_14_), .CO(
        add_6_root_add_0_root_add_94_carry_15_), .S(
        add_6_root_add_0_root_add_94_SUM_14_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_15 ( .A(m27_15_), .B(m29_15_), .CI(
        add_6_root_add_0_root_add_94_carry_15_), .CO(
        add_6_root_add_0_root_add_94_carry_16_), .S(
        add_6_root_add_0_root_add_94_SUM_15_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_16 ( .A(m27_16_), .B(m29_16_), .CI(
        add_6_root_add_0_root_add_94_carry_16_), .CO(
        add_6_root_add_0_root_add_94_carry_17_), .S(
        add_6_root_add_0_root_add_94_SUM_16_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_17 ( .A(m27_17_), .B(m29_17_), .CI(
        add_6_root_add_0_root_add_94_carry_17_), .CO(
        add_6_root_add_0_root_add_94_carry_18_), .S(
        add_6_root_add_0_root_add_94_SUM_17_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_18 ( .A(m27_18_), .B(m29_18_), .CI(
        add_6_root_add_0_root_add_94_carry_18_), .CO(
        add_6_root_add_0_root_add_94_carry_19_), .S(
        add_6_root_add_0_root_add_94_SUM_18_) );
  FA_X1 add_6_root_add_0_root_add_94_U1_19 ( .A(m27_19_), .B(m29_19_), .CI(
        add_6_root_add_0_root_add_94_carry_19_), .CO(
        add_6_root_add_0_root_add_94_carry_20_), .S(
        add_6_root_add_0_root_add_94_SUM_19_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_5 ( .A(m6[2]), .B(m14[1]), .CI(
        add_13_root_add_0_root_add_94_carry[5]), .CO(
        add_13_root_add_0_root_add_94_carry[6]), .S(m29_5_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_6 ( .A(m6[3]), .B(m14[2]), .CI(
        add_13_root_add_0_root_add_94_carry[6]), .CO(
        add_13_root_add_0_root_add_94_carry[7]), .S(m29_6_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_7 ( .A(m6[4]), .B(m14[3]), .CI(
        add_13_root_add_0_root_add_94_carry[7]), .CO(
        add_13_root_add_0_root_add_94_carry[8]), .S(m29_7_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_8 ( .A(m6[5]), .B(m14[4]), .CI(
        add_13_root_add_0_root_add_94_carry[8]), .CO(
        add_13_root_add_0_root_add_94_carry[9]), .S(m29_8_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_9 ( .A(m6[6]), .B(m14[5]), .CI(
        add_13_root_add_0_root_add_94_carry[9]), .CO(
        add_13_root_add_0_root_add_94_carry[10]), .S(m29_9_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_10 ( .A(m6[7]), .B(m14[6]), .CI(
        add_13_root_add_0_root_add_94_carry[10]), .CO(
        add_13_root_add_0_root_add_94_carry[11]), .S(m29_10_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_11 ( .A(m6[8]), .B(m14[7]), .CI(
        add_13_root_add_0_root_add_94_carry[11]), .CO(
        add_13_root_add_0_root_add_94_carry[12]), .S(m29_11_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_12 ( .A(m6[9]), .B(m14[8]), .CI(
        add_13_root_add_0_root_add_94_carry[12]), .CO(
        add_13_root_add_0_root_add_94_carry[13]), .S(m29_12_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_13 ( .A(m6[10]), .B(m14[9]), .CI(
        add_13_root_add_0_root_add_94_carry[13]), .CO(
        add_13_root_add_0_root_add_94_carry[14]), .S(m29_13_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_14 ( .A(m6[11]), .B(m14[10]), .CI(
        add_13_root_add_0_root_add_94_carry[14]), .CO(
        add_13_root_add_0_root_add_94_carry[15]), .S(m29_14_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_15 ( .A(m6[12]), .B(m14[11]), .CI(
        add_13_root_add_0_root_add_94_carry[15]), .CO(
        add_13_root_add_0_root_add_94_carry[16]), .S(m29_15_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_16 ( .A(m6[13]), .B(m14[12]), .CI(
        add_13_root_add_0_root_add_94_carry[16]), .CO(
        add_13_root_add_0_root_add_94_carry[17]), .S(m29_16_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_17 ( .A(m6[14]), .B(m14[13]), .CI(
        add_13_root_add_0_root_add_94_carry[17]), .CO(
        add_13_root_add_0_root_add_94_carry[18]), .S(m29_17_) );
  FA_X1 add_13_root_add_0_root_add_94_U1_18 ( .A(m6[15]), .B(m14[14]), .CI(
        add_13_root_add_0_root_add_94_carry[18]), .CO(
        add_13_root_add_0_root_add_94_carry[19]), .S(m29_18_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_2 ( .A(m18_2_), .B(m24_2_), .CI(
        add_12_root_add_0_root_add_94_carry[2]), .CO(
        add_12_root_add_0_root_add_94_carry[3]), .S(m39_2_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_3 ( .A(m18_3_), .B(m24_3_), .CI(
        add_12_root_add_0_root_add_94_carry[3]), .CO(
        add_12_root_add_0_root_add_94_carry[4]), .S(m39_3_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_4 ( .A(m18_4_), .B(m24_4_), .CI(
        add_12_root_add_0_root_add_94_carry[4]), .CO(
        add_12_root_add_0_root_add_94_carry[5]), .S(m39_4_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_5 ( .A(m18_5_), .B(m24_5_), .CI(
        add_12_root_add_0_root_add_94_carry[5]), .CO(
        add_12_root_add_0_root_add_94_carry[6]), .S(m39_5_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_6 ( .A(m18_6_), .B(m24_6_), .CI(
        add_12_root_add_0_root_add_94_carry[6]), .CO(
        add_12_root_add_0_root_add_94_carry[7]), .S(m39_6_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_7 ( .A(m18_7_), .B(m24_7_), .CI(
        add_12_root_add_0_root_add_94_carry[7]), .CO(
        add_12_root_add_0_root_add_94_carry[8]), .S(m39_7_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_8 ( .A(m18_8_), .B(m24_8_), .CI(
        add_12_root_add_0_root_add_94_carry[8]), .CO(
        add_12_root_add_0_root_add_94_carry[9]), .S(m39_8_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_9 ( .A(m18_9_), .B(m24_9_), .CI(
        add_12_root_add_0_root_add_94_carry[9]), .CO(
        add_12_root_add_0_root_add_94_carry[10]), .S(m39_9_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_10 ( .A(m18_10_), .B(m24_10_), .CI(
        add_12_root_add_0_root_add_94_carry[10]), .CO(
        add_12_root_add_0_root_add_94_carry[11]), .S(m39_10_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_11 ( .A(m18_11_), .B(m24_11_), .CI(
        add_12_root_add_0_root_add_94_carry[11]), .CO(
        add_12_root_add_0_root_add_94_carry[12]), .S(m39_11_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_12 ( .A(m18_12_), .B(m24_12_), .CI(
        add_12_root_add_0_root_add_94_carry[12]), .CO(
        add_12_root_add_0_root_add_94_carry[13]), .S(m39_12_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_13 ( .A(m18_13_), .B(m24_13_), .CI(
        add_12_root_add_0_root_add_94_carry[13]), .CO(
        add_12_root_add_0_root_add_94_carry[14]), .S(m39_13_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_14 ( .A(m18_14_), .B(m24_14_), .CI(
        add_12_root_add_0_root_add_94_carry[14]), .CO(
        add_12_root_add_0_root_add_94_carry[15]), .S(m39_14_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_15 ( .A(m18_15_), .B(m24_15_), .CI(
        add_12_root_add_0_root_add_94_carry[15]), .CO(
        add_12_root_add_0_root_add_94_carry[16]), .S(m39_15_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_16 ( .A(m18_16_), .B(m24_16_), .CI(
        add_12_root_add_0_root_add_94_carry[16]), .CO(
        add_12_root_add_0_root_add_94_carry[17]), .S(m39_16_) );
  FA_X1 add_12_root_add_0_root_add_94_U1_17 ( .A(m18_17_), .B(m24_17_), .CI(
        add_12_root_add_0_root_add_94_carry[17]), .CO(
        add_12_root_add_0_root_add_94_carry[18]), .S(m39_17_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_3 ( .A(m36_3_), .B(m30_3_), .CI(
        add_9_root_add_0_root_add_94_carry[3]), .CO(
        add_9_root_add_0_root_add_94_carry[4]), .S(m37_3_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_4 ( .A(m36_4_), .B(m30_4_), .CI(
        add_9_root_add_0_root_add_94_carry[4]), .CO(
        add_9_root_add_0_root_add_94_carry[5]), .S(m37_4_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_5 ( .A(m36_5_), .B(m30_5_), .CI(
        add_9_root_add_0_root_add_94_carry[5]), .CO(
        add_9_root_add_0_root_add_94_carry[6]), .S(m37_5_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_6 ( .A(m36_6_), .B(m30_6_), .CI(
        add_9_root_add_0_root_add_94_carry[6]), .CO(
        add_9_root_add_0_root_add_94_carry[7]), .S(m37_6_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_7 ( .A(m36_7_), .B(m30_7_), .CI(
        add_9_root_add_0_root_add_94_carry[7]), .CO(
        add_9_root_add_0_root_add_94_carry[8]), .S(m37_7_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_8 ( .A(m36_8_), .B(m30_8_), .CI(
        add_9_root_add_0_root_add_94_carry[8]), .CO(
        add_9_root_add_0_root_add_94_carry[9]), .S(m37_8_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_9 ( .A(m36_9_), .B(m30_9_), .CI(
        add_9_root_add_0_root_add_94_carry[9]), .CO(
        add_9_root_add_0_root_add_94_carry[10]), .S(m37_9_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_10 ( .A(m36_10_), .B(m30_10_), .CI(
        add_9_root_add_0_root_add_94_carry[10]), .CO(
        add_9_root_add_0_root_add_94_carry[11]), .S(m37_10_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_11 ( .A(m36_11_), .B(m30_11_), .CI(
        add_9_root_add_0_root_add_94_carry[11]), .CO(
        add_9_root_add_0_root_add_94_carry[12]), .S(m37_11_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_12 ( .A(m36_12_), .B(m30_12_), .CI(
        add_9_root_add_0_root_add_94_carry[12]), .CO(
        add_9_root_add_0_root_add_94_carry[13]), .S(m37_12_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_13 ( .A(m36_13_), .B(m30_13_), .CI(
        add_9_root_add_0_root_add_94_carry[13]), .CO(
        add_9_root_add_0_root_add_94_carry[14]), .S(m37_13_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_14 ( .A(m36_14_), .B(m30_14_), .CI(
        add_9_root_add_0_root_add_94_carry[14]), .CO(
        add_9_root_add_0_root_add_94_carry[15]), .S(m37_14_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_15 ( .A(m36_15_), .B(m30_15_), .CI(
        add_9_root_add_0_root_add_94_carry[15]), .CO(
        add_9_root_add_0_root_add_94_carry[16]), .S(m37_15_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_16 ( .A(m36_16_), .B(m30_16_), .CI(
        add_9_root_add_0_root_add_94_carry[16]), .CO(
        add_9_root_add_0_root_add_94_carry[17]), .S(m37_16_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_17 ( .A(m36_17_), .B(m30_17_), .CI(
        add_9_root_add_0_root_add_94_carry[17]), .CO(
        add_9_root_add_0_root_add_94_carry[18]), .S(m37_17_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_18 ( .A(m36_18_), .B(m30_18_), .CI(
        add_9_root_add_0_root_add_94_carry[18]), .CO(
        add_9_root_add_0_root_add_94_carry[19]), .S(m37_18_) );
  FA_X1 add_9_root_add_0_root_add_94_U1_19 ( .A(m36_19_), .B(m30_19_), .CI(
        add_9_root_add_0_root_add_94_carry[19]), .CO(m37_20_), .S(m37_19_) );
  INV_X1 U3 ( .A(1'b1), .ZN(y[27]) );
  INV_X1 U5 ( .A(1'b1), .ZN(y[28]) );
  INV_X1 U7 ( .A(1'b1), .ZN(y[29]) );
  INV_X1 U9 ( .A(1'b1), .ZN(y[30]) );
  INV_X1 U11 ( .A(1'b1), .ZN(y[31]) );
  AND2_X1 U13 ( .A1(m42_0_), .A2(m34_0_), .ZN(
        add_8_root_add_0_root_add_94_carry[1]) );
  XOR2_X1 U14 ( .A(m42_0_), .B(m34_0_), .Z(m43_0_) );
  AND2_X1 U15 ( .A1(add_12_root_add_0_root_add_94_carry[18]), .A2(m24_18_), 
        .ZN(m39_19_) );
  XOR2_X1 U16 ( .A(m24_18_), .B(add_12_root_add_0_root_add_94_carry[18]), .Z(
        m39_18_) );
  AND2_X1 U17 ( .A1(m24_1_), .A2(m18_1_), .ZN(
        add_12_root_add_0_root_add_94_carry[2]) );
  XOR2_X1 U18 ( .A(m24_1_), .B(m18_1_), .Z(m39_1_) );
  AND2_X1 U19 ( .A1(m30_2_), .A2(m36_2_), .ZN(
        add_9_root_add_0_root_add_94_carry[3]) );
  XOR2_X1 U20 ( .A(m30_2_), .B(m36_2_), .Z(m37_2_) );
  AND2_X1 U21 ( .A1(add_6_root_add_0_root_add_94_carry_20_), .A2(m29_20_), 
        .ZN(add_6_root_add_0_root_add_94_carry_21_) );
  XOR2_X1 U22 ( .A(m29_20_), .B(add_6_root_add_0_root_add_94_carry_20_), .Z(
        add_6_root_add_0_root_add_94_SUM_20_) );
  AND2_X1 U23 ( .A1(m27_3_), .A2(m29_3_), .ZN(
        add_6_root_add_0_root_add_94_carry_4_) );
  XOR2_X1 U24 ( .A(m29_3_), .B(m27_3_), .Z(add_6_root_add_0_root_add_94_SUM_3_) );
  AND2_X1 U25 ( .A1(add_13_root_add_0_root_add_94_carry[19]), .A2(m14[15]), 
        .ZN(m29_20_) );
  XOR2_X1 U26 ( .A(m14[15]), .B(add_13_root_add_0_root_add_94_carry[19]), .Z(
        m29_19_) );
  AND2_X1 U27 ( .A1(m14[0]), .A2(m6[1]), .ZN(
        add_13_root_add_0_root_add_94_carry[5]) );
  XOR2_X1 U28 ( .A(m14[0]), .B(m6[1]), .Z(m29_4_) );
  AND2_X1 U29 ( .A1(add_14_root_add_0_root_add_94_carry[17]), .A2(m2[15]), 
        .ZN(m31_18_) );
  XOR2_X1 U30 ( .A(m2[15]), .B(add_14_root_add_0_root_add_94_carry[17]), .Z(
        m31_17_) );
  AND2_X1 U31 ( .A1(m2[0]), .A2(m0[1]), .ZN(
        add_14_root_add_0_root_add_94_carry[3]) );
  XOR2_X1 U32 ( .A(m2[0]), .B(m0[1]), .Z(m31_2_) );
endmodule

